module vraphql_enum

pub interface VraphQLEnum {
	value string
}
